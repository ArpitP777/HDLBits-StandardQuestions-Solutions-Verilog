module top_module (
    input clk,
    input slowena,
    input reset,
    output [3:0] q);
    
    always@(posedge clk) begin
        if(reset == 1'b1) begin
            q <= 4'd0;
        end
        else begin
            if(slowena) begin
                if(q == 4'd9)begin
                   q <= 4'd0; 
                end
                else begin
                   q <= q + 4'd1; 
                end
            end
        end
    end

endmodule
